`ifndef INC_PKGS_VH_
    `define INC_PKGS_VH_
    package vproc_pkg;
`endif

